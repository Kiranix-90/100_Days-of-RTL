`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 22.03.2025 19:45:36
// Design Name: 
// Module Name: encoder_8to3
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module encoder_8to3(A7,A6,A5,A4,A3,A2,A1,A0,B,C,D);
input A7,A6,A5,A4,A3,A2,A1,A0;
output B,C,D;

assign B=(A4|A5|A6|A7);
assign C=(A2|A3|A6|A7);
assign D=(A1|A3|A5|A7);

endmodule